���  �A� �                                                �0 ������            �     �                                                 �   �f1����             @     �                                                �   �� ����                   ��                    8       `           p(       � �`  ���                   ��                    l       x           0$       �  �  ����                   �\                    H                   H       � �  �� �                   xt                    4                             `  �� �� ~T                   <                                                  ���� ~             �                                                        �����             �                                       �                �  ���                  �                            p    �                  ���                         �                  �    �             $      ���        �                �                  �� ; -`            ;�    � �        < �      �        �    `             ���x�v             ?��� � � �        @ � � `   �        p1�<�              ��������             �����d� �          < �`              @x����             ��������            ���������                             @����            ���������      �    ���������  <      p                   �   ����           ���������     �    ���������      �       �          �   ~�����          ?���������     �    ?���������� �     �                   �  �����          ��������     �   ���������� �x     a�                 ?�� �?�� `          ` ��������     �   ����������  `|      �                 ?��  �� � �          � �������x     �   ?���������   �     @W�       �          ��  �              � ��������     �   =���������    �     @�                ���      >          �  �������     �   x< ��������  �     ���          @     ����         `     �  }�������   `�   P }������@`p}�     ����      �   �     �����    ��  p     �   y�������  P�   @  y�����������      ���        p0�     ���    ��      �  � ��������� 0  �@   �������������       �        x p  @  ���� ���         � �������`8  �@   �����������  �  � � � �   �   �  ?���   ��      �  �a�����������   �   ��������!����@  @� �      ?�   �  �'��  ��x         �{����������?�   �    �������������       �    ?�      ����  {���   �     ������ ?���/�       �������?��?�0�        {�  ��     ����  s��f         ������ ���=�      ������?�����8�   �   s����     ��?�  G�<  @     ���������� �      <�?����������|�   �   G�< ���     >|��  �8        ��_��������p�     >������������   !��   �8 ��     ?|��    �        ?����������1�    �������� ����    � �     � ��     ����  8 ��         ?�����������    � ��������������   @C     8 � ��     ����  0 �          ���������O���    �����������O�A���    #     0 �        ���� � 	��        �������?�����     p�������?���~" ���        � 	��       ����� � ���        �������?� ��@    �x������?�<����   �2    � ��         ����� ��;��        ������?��?�� d  ��������?�y�?�a���   �!    ��;�  �     ��� ��s��  ��   ����� ��?��� ������ ��?�1��     �!�   �s� �     ���  d����@�   �������?���  ��������?��     �!�    d����     ����  b��O����   �������� 9����  ���������9�����      1�    b`�@ @�     ����  ����  ��   �������  ��� �  ������������      9�    ��  �	�     ����  ��{��  �  �������  ���� ��   �������g�������      9�    �{  7��     �����  ��y�   �  �ۿ�����  ���߀��  @��������������      8�    �y   O�     ���� �����q� �  ������x������  @��?����z������      `@   ��� p�     P_�� ������� �   p_����x<�����   
����x=��_��     ��`   ��� ��     `?�� ǁ����� �   �p����8~  �����    ����8~  �����     ��    ǁ��  �     ��?�� ?����?��� �   �x?���� ~ ��� �   ~������~���_��     ��    >��?  �     ~�?����������� �   �����@  ?�� �   ~����C��?�C��     �   ����<<     >�?����������p �   ~w����    �� �   >�?�������K��     A�   ���~ 4     |�g����������       |g����    ��     <�'�����������   C�x  �G�~d\�   ������������      |�����   � ��      ���'�ǀ�����   #��  �G�8g��   <�����������      =���  0 <� ��    � ����0e������  @#��� G�o ��  `�_���������     �;�����    ?� ��      ����?�t�|�  `��`  � �� ��   ?������������    p���p    ?� �       qо?�|y��   ���/A� ���@�   . ���������    0���0    � �     (   ������   � ��?@���� �   � ������ x~��      |��   ���� �    &�    ���	���|��  x ���  `x ���   �  ����  <<�     <?��   �����x    |0   @��8�����d�   �  ��   < A'��   �  ?���� 0~0    >���   �������    8  `��8����|��   �  {�   >0B�8�   �  ?���� ��0    ~���   ������  �p  a��p������   !�� s�  ~�38�,  �  �����������  3�����   À    ��>`  c0�x3� ��A�� s�  L������@ G�����������ٴ  �����   �   &H  � �   � �hL&h����  � @3����ٔ��  ���������������� � �        d  �0�� ��<��b#D  �� a    �����    ������������������� �       l  ��� �y<�a?� L  ���| a�   �`����    ���������������0�?�� � ��      �  ?��A� ��4����"��  ���x pN  @ �   `	����������������� ?� �>��      L  �@�T� ��<`���`|  �� �0 bN     ���   �������������������=8 '����      L  �@8H@  �`�>��T  ��#Ǉ� �H     �W�    <��� ������������� �1����      \  � ?�@  P@���@  �  �        �?�    8��x ������������� �<����x8�    x  � ?��    < ?��D  � @��        ?�!�    �_��x ������������� ������}��    8  � s�p   "     �E�  � ���        ?� �   ?�a� ?������������ ����������    `0  � �Ā        �f  � -8y�  �      �L�    N� �`=����������`����������    �  � ���        �:�  � }Hx�  �      ��h    ��z 0`=���������� 0���������    �   4x         ����   ɇ�p  B        �d   /��  x���������� ����������    �   �`        ���  	�p            w�   ��� ����������������������    �8����`        ���,  �!��          u������ ?���������Ȝ� �����������    �l����        ���� X  ��� ��          =��A����|��������,���������     x��c��       ����h  ��B� �           ?�� ������<���������$��/p �������     8���7 `       ����$  �����`           /�� ������|���������d���p �������     < �����       �����d  ��o             7�� ������}���������$���� ������     |��� �       ���    ��?             ?�� ?�����?��������� �@� ?������     | ��� q��      ���?$  ��ߎ             �� �����?���������$��� ������    �����@��      ���   �?��     @       �� �����?���������$� � ������    ���� ��       ��   ���             ��������?���������<�  >�����    �������       ?�� <  �~              ��������?���������4�� ������    A���� �        ��  0  ��              ��
������?���������4�(�������   ���  �        ?��  0  v�             �� x��� ?���������4  ]��<�������   �����        ?�� 0  ��8           �� (?��� ���������4  ���<�����?��    ���� �        7��    ���<            �� ���� g���������4  ��~?����'?�    ���(�          ��>0  ��|            ��  ���� ����������4  ��~�����g?�  ���� �         	�~0  ���~           '�� @���� ����������4  �`�������   N��          �0  ��~           �� A���� ����������4  � �~����0��   F�� �         �0  ��~   8        �� �e���� ���������4  ��z�~?���  ��  ���D �         �0  ���~  0        ��D���������������<  8p@���  �  ���t��         � ?�,  ���   p        �� 8�������������<  (�@����   �   >���         | ?�,  ���  �        �� (�����?���������<  � ����       �(�        | ?�(  ���  �        �� A���������������x  @� ����`      ��A��         p�_�l  ��p            �� q��������������x  �q�����`      ��p��         0P�l  ��pAL            ��3?��������������x��1������       �2��        0P?�l����A`            �� #�� �����������x��!� ?�����     0  �"��         ;�L����@            �� �t�� �����������p��#� ;�����      8  ��0ل        �L���� t    @       �� ���� ���������p��� =�����   �p  � !��    @     ������ ~    �      �� ����  ������������� ?�?��   �`  �$ π           ������ ~    �       �� ���  ������������> �� �    �d  ��A��            }�����     �       �� ���  ������������  ?��        l�  À�    �0      <���            �� ���  ������������  ?�?|     � x �  ���     �x      |� ��            �� ���  ?���������� �  ?�?|     �@� �   ��            �|� ~���           �� 	���  ?���������� �  ?� |     0 @� �   ��          �|� {���           �� ����  ?���������� � �� �     �� �  ��             �|� �~���           �� ���   ���������� �`��� �     ��� �  ��            �|���?���            �� ���   ���������� ����� �     ��� �  � 8     �      �|�������           �   ���   �������?�� �`����    �����  �8     �      x�������           �   ��   �������?� ������    ����  ��     �      |��x���           #�   �?p   ?�������?� ��������  @����  ��     �      �����}��           3   �O0   ?�������   �Й�����   ���>   �
�    �      <����=��              ��   �������   ����_���  ���(   � P    �      ������� `           �   �������   ��?���   ���    �;0   � �   ?���w����`            �8��   ?�������   � /���  �?���@   ��y�   �     ?���v�_���         �  �`�   ?�������   ������  �;�#a�F   \���   �     ?���~?���         �  `��   ?������� @� �����  �?�'!�G4  �a��    �     ���p�J���         ��   ���   ?�������   �@� ���  `�o3��$  �('�          _�����?���       ��   ��  �������   � �����  h w�n?c�  �(� 8          �������?���       ��   ��  �������       ����� �x @ ~?A��j%� 8         ����p��?���       �� ���  ��������       ��3��0��   |?R���bPL 8          ���� �,?��        �� ���  ��������      ���c��0��   �����@R �        �����,��         �� '�  ��������     �8���� ��   � 0���Y �        ������&���         �� ��  ��������      �،��� ��  � 0����  �        ����(&���         0����  �� �����      �̏��� ��  � ����P  �        {����,#���         0���~� ��|����      χ�����  ?� ����P �       �?���'����  |     `���>� �� ����     }��������� ����  �        ���~'���� �     ���<� ��|��x     ������.�����N ����8
 (�       1����|���� ��  ���<� ��@   `     {����ǟ������ ����<  8        ��������� ��    ��� � ����        �����ß�<�����   �{�<   ��    �����s���� �      �  x ��opg�      �K��{����p����   ��@ �|  o`    ��������� �g�    �   p ���0�� 8     ����s��� 9����   ��� ��|� �0 #  ��  ���|�� {���� 8   � 0    �� �� 8     ?�������C��   ��� �_�� ` |Ӽ ��  ��~� ����� 8   � �   ������     ��������0��   ��� ;�� ��� ��   ����?� �������   � �   �LX��     �������D�=�   ��� @9� K�X~FB9�`   ����?���������  � �   �?�C����    !������  ?��  ��� �  aC��@?��p   ��������������  �       ������      ���  ��     ��� <�  �����
p   ���?����������  �      �/�����      ����,�     �?�  |� ��J��� �   ������������  �     �82+�����     ���8 (
      ���  |� 82������   ��������������� � �   ��27�����8   ���#��         ��� �` ��2�����'   ���������������� � �   ?������   �?��x  0�     ��� ^�?�����   ����������������� � �   ?��?O���   ���� <<|O�   ���@ � 3�Ã0��   �����������?����� � �  A� ?  ���  ����A� � ǀ ����  =��� 3 �C8x�   ������~��� ������ �  C� ?  � ��   ����
C�  ����     ��  ?�C� 7` �   ��������� � ����� ��  ~  � ��  �����   	���    ��  �  b�� �`�  ����������� � ���� �� $p �`�  x�  �����$p  ��� p   ��  �p 1xv� ���  ��������������� �� �� N   �  ����؁� �Z�<     ��  � � 3� ���  �����?���M ���� �� �0   ��  �����   < �   ��   ��0s@ ��c�  ����������  ���� ����`     xx  �y��� ��d8  `   ��  � h+� ���x  �����c����  � �� ��x@@<       �y���x ��	$ x     ��P &x@ @ۀ ���  ���������<  � �� ����@x��l     �  �}���� ���D <p     ��@ 	�@`  �  ����  ���������|  ���� �?3��?��     �  �}���� ���� 8�  �  �� @3��  (D  ���`  ������?��  �?���  ��d�?�      p  x}�� ���� q� `@  ����d  '   ����  xd����?��  ��|� �����      <   9�� ����0 �� <0  xl�7��   �  ����  =������  ��<� �y�y��         �x ����� �� >  �8�'y�`  
  ���   �������   ��  �������       �  ��� {���w�����  �H-���  �   /���    �������   �?��  �������       �  ߿�����?����d�  � ?��    �    7���    ��������   ���  @w>�W�       �  �w ���߃Ꮐ<�  �  w	�  p  @���    ���?����   ���  A�  ���       �  �� ����#�� > �  � � �   �   ��    ~��?����    ���  C�pp �?�       �  C� 7���g~+�  <    � ��pH  ���   ��    |������    ?� �  Gq�� ��       �  Gp W���gP;�>      ��q��  ���   �   �x�������    ?� � _�À ���       �@_�������|      �8���0 �?�@ ?�   �`?������@     � ��  ��@@      �@������X|      �x?�� �? �  �  ��������     �  ����      �p ��� ��       �x� ���   �  ���� �����     �0�0 1���     � � ���  ��       �z�-� 1��     �  x�� �����     �0�`�  ���     � � @`��  ���       x{�`��� �      �  0��������     � �!� ��       � � � ��  ���       p�!�� �    �  0��������      � �  ��          ����  ���     �0��� �    � � �������         �  ��          �� �� �π     ��_�=�� �    � �  ?�=������         ?�    �@         ?��a�� ��      ����<��     �  ��@�<������        �0    �@          �#�� ��      ��(��      � �����������         �<p    �  @        @� ?����� �\      �~�<@ @     `  `���� �/����        �p�   � �         A� ���� �      �}�p� �    @@     ���� �����        ����             �� ������ ��      �{��  @    @     ���� ������        ���             ���ߟ�� ��      ����  @     @     ��� ������        ᇀ             ������� ��      �/�       �8    ���  ������        �     ��       ������� ��p     �_�     �?��    � ?��  �������       ?�0     �         ?������� �Y�     ���0     �  ���    �@��  �������       p    �0           ������ ���     �`    �  ��    ����|  �������       �0�    �8        �� ������ ���     ��0�    �8 ��� @  ���~  �������       ���   p�,       �� ������� 3���     ���@  @ ���� � @���> @�������       ��   p�`       ��?������ ��      ����    �`��� � @���  ������        �  8p�@@       �������� ?��      ���    �@ �?���  ��� 9������ �      �  8`��A       �������� ?��      ���    �� �?���  ��� 9������ �      ��  8p��A       �����������      ����    � ���   �?��ߜ 9������ @      �8   0p��A       ����������      ��'�    ����  0 ���ߜ 9������            pp A       �  ��������       ��      ��  0 ������ y������        @  Pp       � @��������      �'�      ���$   ������ y������ 8     p�    @p    <   �  ��������   $   �p��    ����   ������ y�������<<     �   @p       � �����������    �� �     ����   ���No� y�������?�     �      p�         � �������� �     �� x    � �����  �� g� y���������     �      p� 	          �������� q       ��    � ����� �  � w��y��������     �     `�           �������� @       ��     @  ���� �  ��w��y�������      �    ` `           ���������`       ��     ` ��� �  ��3��y����=�       �  �  ` @             ������� x       �� �   @ ���� �  � �;�y������                                                                                           ���  �A